module tb_pixel_xformer_avalon();

// Your testbench goes here.

endmodule: tb_pixel_xformer_avalon
