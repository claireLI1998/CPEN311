module tb_task5();

// Your testbench goes here.

endmodule: tb_task5
