module tb_invert_avalon();

// Your testbench goes here.

endmodule: tb_invert_avalon
