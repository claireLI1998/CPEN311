module tb_arc4();

// Your testbench goes here.

endmodule: tb_arc4
