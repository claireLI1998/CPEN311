module tb_prga();

// Your testbench goes here.

endmodule: tb_prga
