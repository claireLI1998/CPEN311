module tb_task4();

// Your testbench goes here.

endmodule: tb_task4
