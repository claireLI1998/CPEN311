module tb_doublecrack();

// Your testbench goes here.

endmodule: tb_doublecrack
