module invert_avalon(input logic clk, input logic reset_n,
                     input logic [3:0] address, input logic write, input logic [31:0] writedata,
                     input logic read, output logic [31:0] readdata);

    // your code here

endmodule: invert_avalon